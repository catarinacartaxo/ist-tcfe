.param V6=7.040227e+00
.param V8=0.0
